LIBRARY ieee;
LIBRARY std;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY ual IS
	GENERIC (N : INTEGER := 32);
	
	PORT (
		
		UALCONTROL : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		SRCA       : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		SRCB       : IN STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		
		RESULT     : OUT STD_LOGIC_VECTOR(N-1 DOWNTO 0);
		COUT       : OUT STD_LOGIC;
		ZERO       : OUT STD_LOGIC
		
	);

END ual;

ARCHITECTURE rtl OF ual IS
	SIGNAL OPERATION : STD_LOGIC_VECTOR(1 DOWNTO 0);
	SIGNAL OP1, OP2  : STD_LOGIC;
	SIGNAL SOMME, SRCA_MUX, SRCB_MUX, RES : STD_LOGIC_VECTOR(N-1 DOWNTO 0);
	SIGNAL RETENUESOMME : UNSIGNED(N DOWNTO 0);
BEGIN

	OPERATION <= UALCONTROL(1 DOWNTO 0);
	OP1       <= UALCONTROL(3);
	OP2       <= UALCONTROL(2);
	
	SRCA_MUX <= NOT(SRCA) WHEN OP1 = '1' ELSE SRCA;
	SRCB_MUX <= NOT(SRCB) WHEN OP2 = '1' ELSE SRCB;
	
	ZERO         <= '1' WHEN SIGNED(RES) = 0 ELSE '0';
	RETENUESOMME <= RESIZE(UNSIGNED(SRCA_MUX), SRCA_MUX'LENGTH+1) + UNSIGNED(SRCB_MUX) + UNSIGNED'("" & OP2);
	SOMME        <= STD_LOGIC_VECTOR(RETENUESOMME(N-1 DOWNTO 0));
	COUT         <= RETENUESOMME(N);
	RESULT       <= RES;
	
	PROCESS (OPERATION, SOMME, SRCA_MUX, SRCB_MUX)
	BEGIN
	
		CASE OPERATION IS
			WHEN "00"   => RES <= STD_LOGIC_VECTOR(SIGNED(SRCA_MUX) AND SIGNED(SRCB_MUX));
			WHEN "01"   => RES <= STD_LOGIC_VECTOR(SIGNED(SRCA_MUX) OR SIGNED(SRCB_MUX));
			WHEN "10"   => RES <= SOMME;
			WHEN "11"   => RES <= (0 => SOMME(N-1), OTHERS => '0');
			WHEN OTHERS => RES <= (OTHERS => 'X');
		END CASE;
	
	END PROCESS;

END RTL;